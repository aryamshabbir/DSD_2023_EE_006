`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/26/2025 10:10:50 PM
// Design Name: 
// Module Name: lab5b
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module lab5b(
  input logic [3:0] num,   
  input logic [2:0] sel,   
  output logic [6:0] segment, 
  output logic [7:0] anode 
    );
 always_comb begin
        case(num)
                4'b0000: segment = 7'b0000001; 
                4'b0001: segment = 7'b1001111; 
                4'b0010: segment = 7'b0010010; 
                4'b0011: segment = 7'b0000110; 
                4'b0100: segment = 7'b1001100; 
                4'b0101: segment = 7'b0100100; 
                4'b0110: segment = 7'b0100000; 
                4'b0111: segment = 7'b0001111; 
                4'b1000: segment = 7'b0000000; 
                4'b1001: segment = 7'b0000100; 
                4'b1010: segment = 7'b0001000; 
                4'b1011: segment = 7'b1100000; 
                4'b1100: segment = 7'b0110001; 
                4'b1101: segment = 7'b1000010; 
                4'b1110: segment = 7'b0110000; 
                4'b1111: segment = 7'b0111000; 
                
          endcase
  end
  always_comb begin
            case(sel)
                3'b000: anode = 8'b11111110; 
                3'b001: anode = 8'b11111101; 
                3'b010: anode = 8'b11111011;
                3'b011: anode = 8'b11110111; 
                3'b100: anode = 8'b11101111; 
                3'b101: anode = 8'b11011111; 
                3'b110: anode = 8'b10111111; 
                3'b111: anode = 8'b01111111; 
                
    endcase
end
        
endmodule
